import ALU::*;

(* synthesize *)
module mkTbALU(Empty);

   function testOne (Bit#(6) fn, Bit#(32) a, Bit#(32) b, Bit#(32) exp) = 
   action
      let got = alu(fn, a, b);
      if (got != exp)
         $display("FAIL fn:%b, a:%h, b:%h, got: %h, expected: %h", fn, a, b, got, exp);
      else
         $display("PASS fn:%b, a:%h, b:%h, got: %h, expected: %h", fn, a, b, got, exp);

   endaction;
   
   rule testAll;
      testOne('b100000, 'hff00ff00, 'hffff0000, 'h00000000);
      testOne('b100001, 'hff00ff00, 'hffff0000, 'h000000ff);
      testOne('b100010, 'hff00ff00, 'hffff0000, 'h0000ff00);
      testOne('b100011, 'hff00ff00, 'hffff0000, 'h0000ffff);
      testOne('b100100, 'hff00ff00, 'hffff0000, 'h00ff0000);
      testOne('b100101, 'hff00ff00, 'hffff0000, 'h00ff00ff);
      testOne('b100110, 'hff00ff00, 'hffff0000, 'h00ffff00);
      testOne('b100111, 'hff00ff00, 'hffff0000, 'h00ffffff);
      testOne('b101000, 'hff00ff00, 'hffff0000, 'hff000000);
      testOne('b101001, 'hff00ff00, 'hffff0000, 'hff0000ff);
      testOne('b101010, 'hff00ff00, 'hffff0000, 'hff00ff00);
      testOne('b101011, 'hff00ff00, 'hffff0000, 'hff00ffff);
      testOne('b101100, 'hff00ff00, 'hffff0000, 'hffff0000);
      testOne('b101101, 'hff00ff00, 'hffff0000, 'hffff00ff);
      testOne('b101110, 'hff00ff00, 'hffff0000, 'hffffff00);
      testOne('b101111, 'hff00ff00, 'hffff0000, 'hffffffff);
      testOne('b110000, 'h00000000, 'h00000000, 'h00000000);
      testOne('b110001, 'h00000000, 'h00000000, 'h00000000);
      testOne('b110011, 'h00000000, 'h00000000, 'h00000000);
      testOne('b110000, 'h00000000, 'h00000001, 'h00000000);
      testOne('b110001, 'h00000000, 'h00000001, 'h00000000);
      testOne('b110011, 'h00000000, 'h00000001, 'h00000000);
      testOne('b110000, 'h00000000, 'h00000002, 'h00000000);
      testOne('b110001, 'h00000000, 'h00000002, 'h00000000);
      testOne('b110011, 'h00000000, 'h00000002, 'h00000000);
      testOne('b110000, 'h00000000, 'h00000004, 'h00000000);
      testOne('b110001, 'h00000000, 'h00000004, 'h00000000);
      testOne('b110011, 'h00000000, 'h00000004, 'h00000000);
      testOne('b110000, 'h00000000, 'h00000008, 'h00000000);
      testOne('b110001, 'h00000000, 'h00000008, 'h00000000);
      testOne('b110011, 'h00000000, 'h00000008, 'h00000000);
      testOne('b110000, 'h00000000, 'h00000010, 'h00000000);
      testOne('b110001, 'h00000000, 'h00000010, 'h00000000);
      testOne('b110011, 'h00000000, 'h00000010, 'h00000000);
      testOne('b110000, 'h00000000, 'h0000001f, 'h00000000);
      testOne('b110001, 'h00000000, 'h0000001f, 'h00000000);
      testOne('b110011, 'h00000000, 'h0000001f, 'h00000000);
      testOne('b110000, 'h00000001, 'h00000000, 'h00000001);
      testOne('b110001, 'h00000001, 'h00000000, 'h00000001);
      testOne('b110011, 'h00000001, 'h00000000, 'h00000001);
      testOne('b110000, 'h00000001, 'h00000001, 'h00000002);
      testOne('b110001, 'h00000001, 'h00000001, 'h00000000);
      testOne('b110011, 'h00000001, 'h00000001, 'h00000000);
      testOne('b110000, 'h00000001, 'h00000002, 'h00000004);
      testOne('b110001, 'h00000001, 'h00000002, 'h00000000);
      testOne('b110011, 'h00000001, 'h00000002, 'h00000000);
      testOne('b110000, 'h00000001, 'h00000004, 'h00000010);
      testOne('b110001, 'h00000001, 'h00000004, 'h00000000);
      testOne('b110011, 'h00000001, 'h00000004, 'h00000000);
      testOne('b110000, 'h00000001, 'h00000008, 'h00000100);
      testOne('b110001, 'h00000001, 'h00000008, 'h00000000);
      testOne('b110011, 'h00000001, 'h00000008, 'h00000000);
      testOne('b110000, 'h00000001, 'h00000010, 'h00010000);
      testOne('b110001, 'h00000001, 'h00000010, 'h00000000);
      testOne('b110011, 'h00000001, 'h00000010, 'h00000000);
      testOne('b110000, 'h00000001, 'h0000001f, 'h80000000);
      testOne('b110001, 'h00000001, 'h0000001f, 'h00000000);
      testOne('b110011, 'h00000001, 'h0000001f, 'h00000000);
      testOne('b110000, 'hffffffff, 'h00000000, 'hffffffff);
      testOne('b110001, 'hffffffff, 'h00000000, 'hffffffff);
      testOne('b110011, 'hffffffff, 'h00000000, 'hffffffff);
      testOne('b110000, 'hffffffff, 'h00000001, 'hfffffffe);
      testOne('b110001, 'hffffffff, 'h00000001, 'h7fffffff);
      testOne('b110011, 'hffffffff, 'h00000001, 'hffffffff);
      testOne('b110000, 'hffffffff, 'h00000002, 'hfffffffc);
      testOne('b110001, 'hffffffff, 'h00000002, 'h3fffffff);
      testOne('b110011, 'hffffffff, 'h00000002, 'hffffffff);
      testOne('b110000, 'hffffffff, 'h00000004, 'hfffffff0);
      testOne('b110001, 'hffffffff, 'h00000004, 'h0fffffff);
      testOne('b110011, 'hffffffff, 'h00000004, 'hffffffff);
      testOne('b110000, 'hffffffff, 'h00000008, 'hffffff00);
      testOne('b110001, 'hffffffff, 'h00000008, 'h00ffffff);
      testOne('b110011, 'hffffffff, 'h00000008, 'hffffffff);
      testOne('b110000, 'hffffffff, 'h00000010, 'hffff0000);
      testOne('b110001, 'hffffffff, 'h00000010, 'h0000ffff);
      testOne('b110011, 'hffffffff, 'h00000010, 'hffffffff);
      testOne('b110000, 'hffffffff, 'h0000001f, 'h80000000);
      testOne('b110001, 'hffffffff, 'h0000001f, 'h00000001);
      testOne('b110011, 'hffffffff, 'h0000001f, 'hffffffff);
      testOne('b110000, 'h12345678, 'h00000000, 'h12345678);
      testOne('b110001, 'h12345678, 'h00000000, 'h12345678);
      testOne('b110011, 'h12345678, 'h00000000, 'h12345678);
      testOne('b110000, 'h12345678, 'h00000001, 'h2468acf0);
      testOne('b110001, 'h12345678, 'h00000001, 'h091a2b3c);
      testOne('b110011, 'h12345678, 'h00000001, 'h091a2b3c);
      testOne('b110000, 'h12345678, 'h00000002, 'h48d159e0);
      testOne('b110001, 'h12345678, 'h00000002, 'h048d159e);
      testOne('b110011, 'h12345678, 'h00000002, 'h048d159e);
      testOne('b110000, 'h12345678, 'h00000004, 'h23456780);
      testOne('b110001, 'h12345678, 'h00000004, 'h01234567);
      testOne('b110011, 'h12345678, 'h00000004, 'h01234567);
      testOne('b110000, 'h12345678, 'h00000008, 'h34567800);
      testOne('b110001, 'h12345678, 'h00000008, 'h00123456);
      testOne('b110011, 'h12345678, 'h00000008, 'h00123456);
      testOne('b110000, 'h12345678, 'h00000010, 'h56780000);
      testOne('b110001, 'h12345678, 'h00000010, 'h00001234);
      testOne('b110011, 'h12345678, 'h00000010, 'h00001234);
      testOne('b110000, 'h12345678, 'h0000001f, 'h00000000);
      testOne('b110001, 'h12345678, 'h0000001f, 'h00000000);
      testOne('b110011, 'h12345678, 'h0000001f, 'h00000000);
      testOne('b110000, 'hfedcab98, 'h00000000, 'hfedcab98);
      testOne('b110001, 'hfedcab98, 'h00000000, 'hfedcab98);
      testOne('b110011, 'hfedcab98, 'h00000000, 'hfedcab98);
      testOne('b110000, 'hfedcab98, 'h00000001, 'hfdb95730);
      testOne('b110001, 'hfedcab98, 'h00000001, 'h7f6e55cc);
      testOne('b110011, 'hfedcab98, 'h00000001, 'hff6e55cc);
      testOne('b110000, 'hfedcab98, 'h00000002, 'hfb72ae60);
      testOne('b110001, 'hfedcab98, 'h00000002, 'h3fb72ae6);
      testOne('b110011, 'hfedcab98, 'h00000002, 'hffb72ae6);
      testOne('b110000, 'hfedcab98, 'h00000004, 'hedcab980);
      testOne('b110001, 'hfedcab98, 'h00000004, 'h0fedcab9);
      testOne('b110011, 'hfedcab98, 'h00000004, 'hffedcab9);
      testOne('b110000, 'hfedcab98, 'h00000008, 'hdcab9800);
      testOne('b110001, 'hfedcab98, 'h00000008, 'h00fedcab);
      testOne('b110011, 'hfedcab98, 'h00000008, 'hfffedcab);
      testOne('b110000, 'hfedcab98, 'h00000010, 'hab980000);
      testOne('b110001, 'hfedcab98, 'h00000010, 'h0000fedc);
      testOne('b110011, 'hfedcab98, 'h00000010, 'hfffffedc);
      testOne('b110000, 'hfedcab98, 'h0000001f, 'h00000000);
      testOne('b110001, 'hfedcab98, 'h0000001f, 'h00000001);
      testOne('b110011, 'hfedcab98, 'h0000001f, 'hffffffff);
      testOne('b010000, 'h00000000, 'h00000000, 'h00000000);
      testOne('b010000, 'h00000000, 'h00000001, 'h00000001);
      testOne('b010000, 'h00000000, 'h-0000001, 'hffffffff);
      testOne('b010000, 'h00000000, 'haaaaaaaa, 'haaaaaaaa);
      testOne('b010000, 'h00000000, 'h55555555, 'h55555555);
      testOne('b010000, 'h00000001, 'h00000000, 'h00000001);
      testOne('b010000, 'h00000001, 'h00000001, 'h00000002);
      testOne('b010000, 'h00000001, 'h-0000001, 'h00000000);
      testOne('b010000, 'h00000001, 'haaaaaaaa, 'haaaaaaab);
      testOne('b010000, 'h00000001, 'h55555555, 'h55555556);
      testOne('b010000, 'h-0000001, 'h00000000, 'hffffffff);
      testOne('b010000, 'h-0000001, 'h00000001, 'h00000000);
      testOne('b010000, 'h-0000001, 'h-0000001, 'hfffffffe);
      testOne('b010000, 'h-0000001, 'haaaaaaaa, 'haaaaaaa9);
      testOne('b010000, 'h-0000001, 'h55555555, 'h55555554);
      testOne('b010000, 'haaaaaaaa, 'h00000000, 'haaaaaaaa);
      testOne('b010000, 'haaaaaaaa, 'h00000001, 'haaaaaaab);
      testOne('b010000, 'haaaaaaaa, 'h-0000001, 'haaaaaaa9);
      testOne('b010000, 'haaaaaaaa, 'haaaaaaaa, 'h55555554);
      testOne('b010000, 'haaaaaaaa, 'h55555555, 'hffffffff);
      testOne('b010000, 'h55555555, 'h00000000, 'h55555555);
      testOne('b010000, 'h55555555, 'h00000001, 'h55555556);
      testOne('b010000, 'h55555555, 'h-0000001, 'h55555554);
      testOne('b010000, 'h55555555, 'haaaaaaaa, 'hffffffff);
      testOne('b010000, 'h55555555, 'h55555555, 'haaaaaaaa);
      testOne('b010001, 'h00000000, 'h00000000, 'h00000000);
      testOne('b010001, 'h00000000, 'h00000001, 'hffffffff);
      testOne('b010001, 'h00000000, 'h-0000001, 'h00000001);
      testOne('b010001, 'h00000000, 'haaaaaaaa, 'h55555556);
      testOne('b010001, 'h00000000, 'h55555555, 'haaaaaaab);
      testOne('b010001, 'h00000001, 'h00000000, 'h00000001);
      testOne('b010001, 'h00000001, 'h00000001, 'h00000000);
      testOne('b010001, 'h00000001, 'h-0000001, 'h00000002);
      testOne('b010001, 'h00000001, 'haaaaaaaa, 'h55555557);
      testOne('b010001, 'h00000001, 'h55555555, 'haaaaaaac);
      testOne('b010001, 'h-0000001, 'h00000000, 'hffffffff);
      testOne('b010001, 'h-0000001, 'h00000001, 'hfffffffe);
      testOne('b010001, 'h-0000001, 'h-0000001, 'h00000000);
      testOne('b010001, 'h-0000001, 'haaaaaaaa, 'h55555555);
      testOne('b010001, 'h-0000001, 'h55555555, 'haaaaaaaa);
      testOne('b010001, 'haaaaaaaa, 'h00000000, 'haaaaaaaa);
      testOne('b010001, 'haaaaaaaa, 'h00000001, 'haaaaaaa9);
      testOne('b010001, 'haaaaaaaa, 'h-0000001, 'haaaaaaab);
      testOne('b010001, 'haaaaaaaa, 'haaaaaaaa, 'h00000000);
      testOne('b010001, 'haaaaaaaa, 'h55555555, 'h55555555);
      testOne('b010001, 'h55555555, 'h00000000, 'h55555555);
      testOne('b010001, 'h55555555, 'h00000001, 'h55555554);
      testOne('b010001, 'h55555555, 'h-0000001, 'h55555556);
      testOne('b010001, 'h55555555, 'haaaaaaaa, 'haaaaaaab);
      testOne('b010001, 'h55555555, 'h55555555, 'h00000000);
      testOne('b000011, 'h00000005, 'hdeadbeef, 'h00000000);
      testOne('b000101, 'h00000005, 'hdeadbeef, 'h00000000);
      testOne('b000111, 'h00000005, 'hdeadbeef, 'h00000000);
      testOne('b000011, 'h12345678, 'h12345678, 'h00000001);
      testOne('b000101, 'h12345678, 'h12345678, 'h00000000);
      testOne('b000111, 'h12345678, 'h12345678, 'h00000001);
      testOne('b000011, 'h80000000, 'h00000001, 'h00000000);
      testOne('b000101, 'h80000000, 'h00000001, 'h00000001);
      testOne('b000111, 'h80000000, 'h00000001, 'h00000001);
      testOne('b000011, 'hdeadbeef, 'h00000005, 'h00000000);
      testOne('b000101, 'hdeadbeef, 'h00000005, 'h00000001);
      testOne('b000111, 'hdeadbeef, 'h00000005, 'h00000001);
      testOne('b000011, 'h7fffffff, 'hffffffff, 'h00000000);
      testOne('b000101, 'h7fffffff, 'hffffffff, 'h00000000);
      testOne('b000111, 'h7fffffff, 'hffffffff, 'h00000000);
      $finish();
   endrule
   
endmodule
