// .power Vdd=1
// .thresholds Vol=0 Vil=0.1 Vih=0.9 Voh=1
// .group inputs SFN[1:0] A[31:0] B[4:0]
// .group outputs Y[31:0]
// .mode gate
// .cycle assert inputs tran 99n sample outputs tran 1n

import Shift::*;

(* synthesize *)
module mkTbShift(Empty);

   function testOne (Bit#(2) sfn, Bit#(32) a, Bit#(5) b, Bit#(32) exp) = 
   action
      let got = shift(sfn, a, b);
      if (got != exp)
         $display("FAIL sfn:%b, a:%b, b:%b, got: %b, expected: %b", sfn, a, b, got, exp);
      else
         $display("PASS sfn:%b, a:%b, b:%b, got: %b, expected: %b", sfn, a, b, got, exp);
   endaction;

   rule testAll;
      testOne('b00, 'h00000000, 'b00000, 'h00000000);
      testOne('b01, 'h00000000, 'b00000, 'h00000000);
      testOne('b11, 'h00000000, 'b00000, 'h00000000);
      testOne('b00, 'h00000000, 'b00001, 'h00000000);
      testOne('b01, 'h00000000, 'b00001, 'h00000000);
      testOne('b11, 'h00000000, 'b00001, 'h00000000);
      testOne('b00, 'h00000000, 'b00010, 'h00000000);
      testOne('b01, 'h00000000, 'b00010, 'h00000000);
      testOne('b11, 'h00000000, 'b00010, 'h00000000);
      testOne('b00, 'h00000000, 'b00100, 'h00000000);
      testOne('b01, 'h00000000, 'b00100, 'h00000000);
      testOne('b11, 'h00000000, 'b00100, 'h00000000);
      testOne('b00, 'h00000000, 'b01000, 'h00000000);
      testOne('b01, 'h00000000, 'b01000, 'h00000000);
      testOne('b11, 'h00000000, 'b01000, 'h00000000);
      testOne('b00, 'h00000000, 'b10000, 'h00000000);
      testOne('b01, 'h00000000, 'b10000, 'h00000000);
      testOne('b11, 'h00000000, 'b10000, 'h00000000);
      testOne('b00, 'h00000000, 'b11111, 'h00000000);
      testOne('b01, 'h00000000, 'b11111, 'h00000000);
      testOne('b11, 'h00000000, 'b11111, 'h00000000);
      testOne('b00, 'h00000001, 'b00000, 'h00000001);
      testOne('b01, 'h00000001, 'b00000, 'h00000001);
      testOne('b11, 'h00000001, 'b00000, 'h00000001);
      testOne('b00, 'h00000001, 'b00001, 'h00000002);
      testOne('b01, 'h00000001, 'b00001, 'h00000000);
      testOne('b11, 'h00000001, 'b00001, 'h00000000);
      testOne('b00, 'h00000001, 'b00010, 'h00000004);
      testOne('b01, 'h00000001, 'b00010, 'h00000000);
      testOne('b11, 'h00000001, 'b00010, 'h00000000);
      testOne('b00, 'h00000001, 'b00100, 'h00000010);
      testOne('b01, 'h00000001, 'b00100, 'h00000000);
      testOne('b11, 'h00000001, 'b00100, 'h00000000);
      testOne('b00, 'h00000001, 'b01000, 'h00000100);
      testOne('b01, 'h00000001, 'b01000, 'h00000000);
      testOne('b11, 'h00000001, 'b01000, 'h00000000);
      testOne('b00, 'h00000001, 'b10000, 'h00010000);
      testOne('b01, 'h00000001, 'b10000, 'h00000000);
      testOne('b11, 'h00000001, 'b10000, 'h00000000);
      testOne('b00, 'h00000001, 'b11111, 'h80000000);
      testOne('b01, 'h00000001, 'b11111, 'h00000000);
      testOne('b11, 'h00000001, 'b11111, 'h00000000);
      testOne('b00, 'hFFFFFFFF, 'b00000, 'hFFFFFFFF);
      testOne('b01, 'hFFFFFFFF, 'b00000, 'hFFFFFFFF);
      testOne('b11, 'hFFFFFFFF, 'b00000, 'hFFFFFFFF);
      testOne('b00, 'hFFFFFFFF, 'b00001, 'hFFFFFFFE);
      testOne('b01, 'hFFFFFFFF, 'b00001, 'h7FFFFFFF);
      testOne('b11, 'hFFFFFFFF, 'b00001, 'hFFFFFFFF);
      testOne('b00, 'hFFFFFFFF, 'b00010, 'hFFFFFFFC);
      testOne('b01, 'hFFFFFFFF, 'b00010, 'h3FFFFFFF);
      testOne('b11, 'hFFFFFFFF, 'b00010, 'hFFFFFFFF);
      testOne('b00, 'hFFFFFFFF, 'b00100, 'hFFFFFFF0);
      testOne('b01, 'hFFFFFFFF, 'b00100, 'h0FFFFFFF);
      testOne('b11, 'hFFFFFFFF, 'b00100, 'hFFFFFFFF);
      testOne('b00, 'hFFFFFFFF, 'b01000, 'hFFFFFF00);
      testOne('b01, 'hFFFFFFFF, 'b01000, 'h00FFFFFF);
      testOne('b11, 'hFFFFFFFF, 'b01000, 'hFFFFFFFF);
      testOne('b00, 'hFFFFFFFF, 'b10000, 'hFFFF0000);
      testOne('b01, 'hFFFFFFFF, 'b10000, 'h0000FFFF);
      testOne('b11, 'hFFFFFFFF, 'b10000, 'hFFFFFFFF);
      testOne('b00, 'hFFFFFFFF, 'b11111, 'h80000000);
      testOne('b01, 'hFFFFFFFF, 'b11111, 'h00000001);
      testOne('b11, 'hFFFFFFFF, 'b11111, 'hFFFFFFFF);
      testOne('b00, 'h12345678, 'b00000, 'h12345678);
      testOne('b01, 'h12345678, 'b00000, 'h12345678);
      testOne('b11, 'h12345678, 'b00000, 'h12345678);
      testOne('b00, 'h12345678, 'b00001, 'h2468ACF0);
      testOne('b01, 'h12345678, 'b00001, 'h091A2B3C);
      testOne('b11, 'h12345678, 'b00001, 'h091A2B3C);
      testOne('b00, 'h12345678, 'b00010, 'h48D159E0);
      testOne('b01, 'h12345678, 'b00010, 'h048D159E);
      testOne('b11, 'h12345678, 'b00010, 'h048D159E);
      testOne('b00, 'h12345678, 'b00100, 'h23456780);
      testOne('b01, 'h12345678, 'b00100, 'h01234567);
      testOne('b11, 'h12345678, 'b00100, 'h01234567);
      testOne('b00, 'h12345678, 'b01000, 'h34567800);
      testOne('b01, 'h12345678, 'b01000, 'h00123456);
      testOne('b11, 'h12345678, 'b01000, 'h00123456);
      testOne('b00, 'h12345678, 'b10000, 'h56780000);
      testOne('b01, 'h12345678, 'b10000, 'h00001234);
      testOne('b11, 'h12345678, 'b10000, 'h00001234);
      testOne('b00, 'h12345678, 'b11111, 'h00000000);
      testOne('b01, 'h12345678, 'b11111, 'h00000000);
      testOne('b11, 'h12345678, 'b11111, 'h00000000);
      testOne('b00, 'hFEDCBA98, 'b00000, 'hFEDCBA98);
      testOne('b01, 'hFEDCBA98, 'b00000, 'hFEDCBA98);
      testOne('b11, 'hFEDCBA98, 'b00000, 'hFEDCBA98);
      testOne('b00, 'hFEDCBA98, 'b00001, 'hFDB97530);
      testOne('b01, 'hFEDCBA98, 'b00001, 'h7F6E5D4C);
      testOne('b11, 'hFEDCBA98, 'b00001, 'hFF6E5D4C);
      testOne('b00, 'hFEDCBA98, 'b00010, 'hFB72EA60);
      testOne('b01, 'hFEDCBA98, 'b00010, 'h3FB72EA6);
      testOne('b11, 'hFEDCBA98, 'b00010, 'hFFB72EA6);
      testOne('b00, 'hFEDCBA98, 'b00100, 'hEDCBA980);
      testOne('b01, 'hFEDCBA98, 'b00100, 'h0FEDCBA9);
      testOne('b11, 'hFEDCBA98, 'b00100, 'hFFEDCBA9);
      testOne('b00, 'hFEDCBA98, 'b01000, 'hDCBA9800);
      testOne('b01, 'hFEDCBA98, 'b01000, 'h00FEDCBA);
      testOne('b11, 'hFEDCBA98, 'b01000, 'hFFFEDCBA);
      testOne('b00, 'hFEDCBA98, 'b10000, 'hBA980000);
      testOne('b01, 'hFEDCBA98, 'b10000, 'h0000FEDC);
      testOne('b11, 'hFEDCBA98, 'b10000, 'hFFFFFEDC);
      testOne('b00, 'hFEDCBA98, 'b11111, 'h00000000);
      testOne('b01, 'hFEDCBA98, 'b11111, 'h00000001);
      testOne('b11, 'hFEDCBA98, 'b11111, 'hFFFFFFFF);
      

      
      $finish();
   endrule
endmodule


// 00 00000000000000000000000000000000 00000 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //   1: fn=SHL, a=0X00000000, b= 0, y=0X00000000
// 01 00000000000000000000000000000000 00000 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //   2: fn=SHR, a=0X00000000, b= 0, y=0X00000000
// 11 00000000000000000000000000000000 00000 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //   3: fn=SRA, a=0X00000000, b= 0, y=0X00000000
// 00 00000000000000000000000000000000 00001 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //   4: fn=SHL, a=0X00000000, b= 1, y=0X00000000
// 01 00000000000000000000000000000000 00001 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //   5: fn=SHR, a=0X00000000, b= 1, y=0X00000000
// 11 00000000000000000000000000000000 00001 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //   6: fn=SRA, a=0X00000000, b= 1, y=0X00000000
// 00 00000000000000000000000000000000 00010 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //   7: fn=SHL, a=0X00000000, b= 2, y=0X00000000
// 01 00000000000000000000000000000000 00010 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //   8: fn=SHR, a=0X00000000, b= 2, y=0X00000000
// 11 00000000000000000000000000000000 00010 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //   9: fn=SRA, a=0X00000000, b= 2, y=0X00000000
// 00 00000000000000000000000000000000 00100 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  10: fn=SHL, a=0X00000000, b= 4, y=0X00000000
// 01 00000000000000000000000000000000 00100 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  11: fn=SHR, a=0X00000000, b= 4, y=0X00000000
// 11 00000000000000000000000000000000 00100 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  12: fn=SRA, a=0X00000000, b= 4, y=0X00000000
// 00 00000000000000000000000000000000 01000 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  13: fn=SHL, a=0X00000000, b= 8, y=0X00000000
// 01 00000000000000000000000000000000 01000 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  14: fn=SHR, a=0X00000000, b= 8, y=0X00000000
// 11 00000000000000000000000000000000 01000 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  15: fn=SRA, a=0X00000000, b= 8, y=0X00000000
// 00 00000000000000000000000000000000 10000 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  16: fn=SHL, a=0X00000000, b=16, y=0X00000000
// 01 00000000000000000000000000000000 10000 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  17: fn=SHR, a=0X00000000, b=16, y=0X00000000
// 11 00000000000000000000000000000000 10000 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  18: fn=SRA, a=0X00000000, b=16, y=0X00000000
// 00 00000000000000000000000000000000 11111 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  19: fn=SHL, a=0X00000000, b=31, y=0X00000000
// 01 00000000000000000000000000000000 11111 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  20: fn=SHR, a=0X00000000, b=31, y=0X00000000
// 11 00000000000000000000000000000000 11111 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  21: fn=SRA, a=0X00000000, b=31, y=0X00000000
// 00 00000000000000000000000000000001 00000 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLH //  22: fn=SHL, a=0X00000001, b= 0, y=0X00000001
// 01 00000000000000000000000000000001 00000 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLH //  23: fn=SHR, a=0X00000001, b= 0, y=0X00000001
// 11 00000000000000000000000000000001 00000 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLH //  24: fn=SRA, a=0X00000001, b= 0, y=0X00000001
// 00 00000000000000000000000000000001 00001 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLHL //  25: fn=SHL, a=0X00000001, b= 1, y=0X00000002
// 01 00000000000000000000000000000001 00001 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  26: fn=SHR, a=0X00000001, b= 1, y=0X00000000
// 11 00000000000000000000000000000001 00001 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  27: fn=SRA, a=0X00000001, b= 1, y=0X00000000
// 00 00000000000000000000000000000001 00010 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLHLL //  28: fn=SHL, a=0X00000001, b= 2, y=0X00000004
// 01 00000000000000000000000000000001 00010 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  29: fn=SHR, a=0X00000001, b= 2, y=0X00000000
// 11 00000000000000000000000000000001 00010 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  30: fn=SRA, a=0X00000001, b= 2, y=0X00000000
// 00 00000000000000000000000000000001 00100 LLLLLLLLLLLLLLLLLLLLLLLLLLLHLLLL //  31: fn=SHL, a=0X00000001, b= 4, y=0X00000010
// 01 00000000000000000000000000000001 00100 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  32: fn=SHR, a=0X00000001, b= 4, y=0X00000000
// 11 00000000000000000000000000000001 00100 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  33: fn=SRA, a=0X00000001, b= 4, y=0X00000000
// 00 00000000000000000000000000000001 01000 LLLLLLLLLLLLLLLLLLLLLLLHLLLLLLLL //  34: fn=SHL, a=0X00000001, b= 8, y=0X00000100
// 01 00000000000000000000000000000001 01000 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  35: fn=SHR, a=0X00000001, b= 8, y=0X00000000
// 11 00000000000000000000000000000001 01000 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  36: fn=SRA, a=0X00000001, b= 8, y=0X00000000
// 00 00000000000000000000000000000001 10000 LLLLLLLLLLLLLLLHLLLLLLLLLLLLLLLL //  37: fn=SHL, a=0X00000001, b=16, y=0X00010000
// 01 00000000000000000000000000000001 10000 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  38: fn=SHR, a=0X00000001, b=16, y=0X00000000
// 11 00000000000000000000000000000001 10000 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  39: fn=SRA, a=0X00000001, b=16, y=0X00000000
// 00 00000000000000000000000000000001 11111 HLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  40: fn=SHL, a=0X00000001, b=31, y=0X80000000
// 01 00000000000000000000000000000001 11111 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  41: fn=SHR, a=0X00000001, b=31, y=0X00000000
// 11 00000000000000000000000000000001 11111 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  42: fn=SRA, a=0X00000001, b=31, y=0X00000000
// 00 11111111111111111111111111111111 00000 HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH //  43: fn=SHL, a=0XFFFFFFFF, b= 0, y=0XFFFFFFFF
// 01 11111111111111111111111111111111 00000 HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH //  44: fn=SHR, a=0XFFFFFFFF, b= 0, y=0XFFFFFFFF
// 11 11111111111111111111111111111111 00000 HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH //  45: fn=SRA, a=0XFFFFFFFF, b= 0, y=0XFFFFFFFF
// 00 11111111111111111111111111111111 00001 HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHL //  46: fn=SHL, a=0XFFFFFFFF, b= 1, y=0XFFFFFFFE
// 01 11111111111111111111111111111111 00001 LHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH //  47: fn=SHR, a=0XFFFFFFFF, b= 1, y=0X7FFFFFFF
// 11 11111111111111111111111111111111 00001 HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH //  48: fn=SRA, a=0XFFFFFFFF, b= 1, y=0XFFFFFFFF
// 00 11111111111111111111111111111111 00010 HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHLL //  49: fn=SHL, a=0XFFFFFFFF, b= 2, y=0XFFFFFFFC
// 01 11111111111111111111111111111111 00010 LLHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH //  50: fn=SHR, a=0XFFFFFFFF, b= 2, y=0X3FFFFFFF
// 11 11111111111111111111111111111111 00010 HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH //  51: fn=SRA, a=0XFFFFFFFF, b= 2, y=0XFFFFFFFF
// 00 11111111111111111111111111111111 00100 HHHHHHHHHHHHHHHHHHHHHHHHHHHHLLLL //  52: fn=SHL, a=0XFFFFFFFF, b= 4, y=0XFFFFFFF0
// 01 11111111111111111111111111111111 00100 LLLLHHHHHHHHHHHHHHHHHHHHHHHHHHHH //  53: fn=SHR, a=0XFFFFFFFF, b= 4, y=0X0FFFFFFF
// 11 11111111111111111111111111111111 00100 HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH //  54: fn=SRA, a=0XFFFFFFFF, b= 4, y=0XFFFFFFFF
// 00 11111111111111111111111111111111 01000 HHHHHHHHHHHHHHHHHHHHHHHHLLLLLLLL //  55: fn=SHL, a=0XFFFFFFFF, b= 8, y=0XFFFFFF00
// 01 11111111111111111111111111111111 01000 LLLLLLLLHHHHHHHHHHHHHHHHHHHHHHHH //  56: fn=SHR, a=0XFFFFFFFF, b= 8, y=0X00FFFFFF
// 11 11111111111111111111111111111111 01000 HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH //  57: fn=SRA, a=0XFFFFFFFF, b= 8, y=0XFFFFFFFF
// 00 11111111111111111111111111111111 10000 HHHHHHHHHHHHHHHHLLLLLLLLLLLLLLLL //  58: fn=SHL, a=0XFFFFFFFF, b=16, y=0XFFFF0000
// 01 11111111111111111111111111111111 10000 LLLLLLLLLLLLLLLLHHHHHHHHHHHHHHHH //  59: fn=SHR, a=0XFFFFFFFF, b=16, y=0X0000FFFF
// 11 11111111111111111111111111111111 10000 HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH //  60: fn=SRA, a=0XFFFFFFFF, b=16, y=0XFFFFFFFF
// 00 11111111111111111111111111111111 11111 HLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  61: fn=SHL, a=0XFFFFFFFF, b=31, y=0X80000000
// 01 11111111111111111111111111111111 11111 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLH //  62: fn=SHR, a=0XFFFFFFFF, b=31, y=0X00000001
// 11 11111111111111111111111111111111 11111 HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH //  63: fn=SRA, a=0XFFFFFFFF, b=31, y=0XFFFFFFFF
// 00 00010010001101000101011001111000 00000 LLLHLLHLLLHHLHLLLHLHLHHLLHHHHLLL //  64: fn=SHL, a=0X12345678, b= 0, y=0X12345678
// 01 00010010001101000101011001111000 00000 LLLHLLHLLLHHLHLLLHLHLHHLLHHHHLLL //  65: fn=SHR, a=0X12345678, b= 0, y=0X12345678
// 11 00010010001101000101011001111000 00000 LLLHLLHLLLHHLHLLLHLHLHHLLHHHHLLL //  66: fn=SRA, a=0X12345678, b= 0, y=0X12345678
// 00 00010010001101000101011001111000 00001 LLHLLHLLLHHLHLLLHLHLHHLLHHHHLLLL //  67: fn=SHL, a=0X12345678, b= 1, y=0X2468ACF0
// 01 00010010001101000101011001111000 00001 LLLLHLLHLLLHHLHLLLHLHLHHLLHHHHLL //  68: fn=SHR, a=0X12345678, b= 1, y=0X091A2B3C
// 11 00010010001101000101011001111000 00001 LLLLHLLHLLLHHLHLLLHLHLHHLLHHHHLL //  69: fn=SRA, a=0X12345678, b= 1, y=0X091A2B3C
// 00 00010010001101000101011001111000 00010 LHLLHLLLHHLHLLLHLHLHHLLHHHHLLLLL //  70: fn=SHL, a=0X12345678, b= 2, y=0X48D159E0
// 01 00010010001101000101011001111000 00010 LLLLLHLLHLLLHHLHLLLHLHLHHLLHHHHL //  71: fn=SHR, a=0X12345678, b= 2, y=0X048D159E
// 11 00010010001101000101011001111000 00010 LLLLLHLLHLLLHHLHLLLHLHLHHLLHHHHL //  72: fn=SRA, a=0X12345678, b= 2, y=0X048D159E
// 00 00010010001101000101011001111000 00100 LLHLLLHHLHLLLHLHLHHLLHHHHLLLLLLL //  73: fn=SHL, a=0X12345678, b= 4, y=0X23456780
// 01 00010010001101000101011001111000 00100 LLLLLLLHLLHLLLHHLHLLLHLHLHHLLHHH //  74: fn=SHR, a=0X12345678, b= 4, y=0X01234567
// 11 00010010001101000101011001111000 00100 LLLLLLLHLLHLLLHHLHLLLHLHLHHLLHHH //  75: fn=SRA, a=0X12345678, b= 4, y=0X01234567
// 00 00010010001101000101011001111000 01000 LLHHLHLLLHLHLHHLLHHHHLLLLLLLLLLL //  76: fn=SHL, a=0X12345678, b= 8, y=0X34567800
// 01 00010010001101000101011001111000 01000 LLLLLLLLLLLHLLHLLLHHLHLLLHLHLHHL //  77: fn=SHR, a=0X12345678, b= 8, y=0X00123456
// 11 00010010001101000101011001111000 01000 LLLLLLLLLLLHLLHLLLHHLHLLLHLHLHHL //  78: fn=SRA, a=0X12345678, b= 8, y=0X00123456
// 00 00010010001101000101011001111000 10000 LHLHLHHLLHHHHLLLLLLLLLLLLLLLLLLL //  79: fn=SHL, a=0X12345678, b=16, y=0X56780000
// 01 00010010001101000101011001111000 10000 LLLLLLLLLLLLLLLLLLLHLLHLLLHHLHLL //  80: fn=SHR, a=0X12345678, b=16, y=0X00001234
// 11 00010010001101000101011001111000 10000 LLLLLLLLLLLLLLLLLLLHLLHLLLHHLHLL //  81: fn=SRA, a=0X12345678, b=16, y=0X00001234
// 00 00010010001101000101011001111000 11111 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  82: fn=SHL, a=0X12345678, b=31, y=0X00000000
// 01 00010010001101000101011001111000 11111 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  83: fn=SHR, a=0X12345678, b=31, y=0X00000000
// 11 00010010001101000101011001111000 11111 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL //  84: fn=SRA, a=0X12345678, b=31, y=0X00000000
// 00 11111110110111001011101010011000 00000 HHHHHHHLHHLHHHLLHLHHHLHLHLLHHLLL //  85: fn=SHL, a=0XFEDCBA98, b= 0, y=0XFEDCBA98
// 01 11111110110111001011101010011000 00000 HHHHHHHLHHLHHHLLHLHHHLHLHLLHHLLL //  86: fn=SHR, a=0XFEDCBA98, b= 0, y=0XFEDCBA98
// 11 11111110110111001011101010011000 00000 HHHHHHHLHHLHHHLLHLHHHLHLHLLHHLLL //  87: fn=SRA, a=0XFEDCBA98, b= 0, y=0XFEDCBA98
// 00 11111110110111001011101010011000 00001 HHHHHHLHHLHHHLLHLHHHLHLHLLHHLLLL //  88: fn=SHL, a=0XFEDCBA98, b= 1, y=0XFDB97530
// 01 11111110110111001011101010011000 00001 LHHHHHHHLHHLHHHLLHLHHHLHLHLLHHLL //  89: fn=SHR, a=0XFEDCBA98, b= 1, y=0X7F6E5D4C
// 11 11111110110111001011101010011000 00001 HHHHHHHHLHHLHHHLLHLHHHLHLHLLHHLL //  90: fn=SRA, a=0XFEDCBA98, b= 1, y=0XFF6E5D4C
// 00 11111110110111001011101010011000 00010 HHHHHLHHLHHHLLHLHHHLHLHLLHHLLLLL //  91: fn=SHL, a=0XFEDCBA98, b= 2, y=0XFB72EA60
// 01 11111110110111001011101010011000 00010 LLHHHHHHHLHHLHHHLLHLHHHLHLHLLHHL //  92: fn=SHR, a=0XFEDCBA98, b= 2, y=0X3FB72EA6
// 11 11111110110111001011101010011000 00010 HHHHHHHHHLHHLHHHLLHLHHHLHLHLLHHL //  93: fn=SRA, a=0XFEDCBA98, b= 2, y=0XFFB72EA6
// 00 11111110110111001011101010011000 00100 HHHLHHLHHHLLHLHHHLHLHLLHHLLLLLLL //  94: fn=SHL, a=0XFEDCBA98, b= 4, y=0XEDCBA980
// 01 11111110110111001011101010011000 00100 LLLLHHHHHHHLHHLHHHLLHLHHHLHLHLLH //  95: fn=SHR, a=0XFEDCBA98, b= 4, y=0X0FEDCBA9
// 11 11111110110111001011101010011000 00100 HHHHHHHHHHHLHHLHHHLLHLHHHLHLHLLH //  96: fn=SRA, a=0XFEDCBA98, b= 4, y=0XFFEDCBA9
// 00 11111110110111001011101010011000 01000 HHLHHHLLHLHHHLHLHLLHHLLLLLLLLLLL //  97: fn=SHL, a=0XFEDCBA98, b= 8, y=0XDCBA9800
// 01 11111110110111001011101010011000 01000 LLLLLLLLHHHHHHHLHHLHHHLLHLHHHLHL //  98: fn=SHR, a=0XFEDCBA98, b= 8, y=0X00FEDCBA
// 11 11111110110111001011101010011000 01000 HHHHHHHHHHHHHHHLHHLHHHLLHLHHHLHL //  99: fn=SRA, a=0XFEDCBA98, b= 8, y=0XFFFEDCBA
// 00 11111110110111001011101010011000 10000 HLHHHLHLHLLHHLLLLLLLLLLLLLLLLLLL // 100: fn=SHL, a=0XFEDCBA98, b=16, y=0XBA980000
// 01 11111110110111001011101010011000 10000 LLLLLLLLLLLLLLLLHHHHHHHLHHLHHHLL // 101: fn=SHR, a=0XFEDCBA98, b=16, y=0X0000FEDC
// 11 11111110110111001011101010011000 10000 HHHHHHHHHHHHHHHHHHHHHHHLHHLHHHLL // 102: fn=SRA, a=0XFEDCBA98, b=16, y=0XFFFFFEDC
// 00 11111110110111001011101010011000 11111 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLL // 103: fn=SHL, a=0XFEDCBA98, b=31, y=0X00000000
// 01 11111110110111001011101010011000 11111 LLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLH // 104: fn=SHR, a=0XFEDCBA98, b=31, y=0X00000001
// 11 11111110110111001011101010011000 11111 HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH // 105: fn=SRA, a=0XFEDCBA98, b=31, y=0XFFFFFFFF
