../Bool.bsv