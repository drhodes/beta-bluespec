import Pc::*;

(* synthesize *)
module mkTbPc(Empty);
   let pcUnit <- mkPc();
   Reg#(Int#(32)) cycle <- mkReg(0);
   
   function testOne(Bit#(1) reset, 
                    Bit#(3) pc_sel, 
                    Bit#(16) id, 
                    Bit#(32) jt, 
                    Bit#(32) pc, 
                    Bit#(32) pc_inc, 
                    Bit#(32) pc_offset) = 
   action
      $display("---- cycle: %d", cycle);
      pcUnit.next(reset, pc_sel, id, jt);
      let result = pcUnit.read(); 
      if (result.pc != pc) begin
         // || result.pc_inc != pc_inc || result.pc_offset != pc_offset) begin
         $display("FAIL reset:%b", reset);
         $display("FAIL pc_sel:%b", pc_sel);
         $display("FAIL id:%h", id);
         $display("FAIL jt:%h", jt);
         $display("FAIL pc:        got: %h, exp: %h", result.pc, pc);
         $display("FAIL pc_inc:    got: %h, exp: %h", result.pc_inc, pc_inc);
         $display("FAIL pc_offset: got: %h, exp: %h", result.pc_offset, pc_offset);
      end
      else $display("PASS pc: got: %h, exp: %h", result.pc, pc);
      cycle <= cycle + 1;
   endaction;
   
   rule t0(cycle == 0);
      $display("resetting unit");
      pcUnit.reset_unit();      
      cycle <= cycle + 1;
   endrule
   
   rule t1(cycle == 1);      
      testOne('b1, 'b011, 'b1111111111111111, 'b00000000000000000000000000000000,
              'b10000000000000000000000000000000,
              'b10000000000000000000000000000100,
              'b10000000000000000000000000000000); //   1: reset, PC==0x80000000
   endrule   
   rule t2(cycle == 2);
      testOne('b1, 'b011, 'b1111111111111111, 'b00000000000000000000000000000000,
              'b10000000000000000000000000000000,
              'b10000000000000000000000000000100,
              'b10000000000000000000000000000000); //   2: reset, PC==0x80000000
   endrule
   rule t3 (cycle == 3);
      testOne('b1, 'b100, 'b0000000000000000, 'b00000000000000000000000000000000,
              'b10000000000000000000000000000000,
              'b10000000000000000000000000000100,
              'b10000000000000000000000000000100); //   3: reset, PC==0x80000000
   endrule
   rule t4 (cycle == 4);
      testOne('b0, 'b100, 'b1111111111111110, 'b00000000000000000000000000000000,
              'b10000000000000000000000000001000,
              'b10000000000000000000000000001100,
              'b10000000000000000000000000000100); //   4: xadr, PC==0x80000008, offset=-2
      $finish();
   endrule
   // rule t5 (cycle == 5);
   //    testOne('b0, 'b011, 'b0111111111111111, 'b00000000000000000000000000000000,
   //            'b10000000000000000000000000000100,
   //            'b10000000000000000000000000001000,
   //            'b10000000000000100000000000000100); //   5: illop, PC==0x80000004, offset=0x7fff
   // endrule
   // rule t6 (cycle == 6);
   //    testOne('b0, 'b010, 'b0000000000000000, 'b11111111111111111111111111110000,
   //            'b11111111111111111111111111110000,
   //            'b11111111111111111111111111110100,
   //            'b11111111111111111111111111110100); //   6: jmp, pc==0XFFFFFFF0
   // endrule
   // rule t7 (cycle == 7);
   //    testOne('b0, 'b000, 'b1111111111111111, 'b00000000000000000000000000000000,
   //            'b11111111111111111111111111110100,
   //            'b11111111111111111111111111111000,
   //            'b11111111111111111111111111110100); //   7: inc, pc==0xFFFFFFF4, offset=-1
   // endrule
   // rule t8 (cycle == 8);
   //    testOne('b0, 'b000, 'b1111111111111110, 'b00000000000000000000000000000000,
   //            'b11111111111111111111111111111000,
   //            'b11111111111111111111111111111100,
   //            'b11111111111111111111111111110100); //   8: inc, pc==0xFFFFFFF8, offset=-1
   // endrule
   // rule t9 (cycle == 9);
   //    testOne('b0, 'b000, 'b1111111111111101, 'b00000000000000000000000000000000,
   //            'b11111111111111111111111111111100,
   //            'b10000000000000000000000000000000,
   //            'b11111111111111111111111111110100); //   9: inc, pc==0xFFFFFFFC, offset=-1
   // endrule
   // rule t10 (cycle == 10);
   //    testOne('b0, 'b000, 'b1111111111111100, 'b00000000000000000000000000000000,
   //            'b10000000000000000000000000000000,
   //            'b10000000000000000000000000000100,
   //            'b11111111111111111111111111110100); //  10: inc, pc==0x80000000, offset=-1
   // endrule
   // rule t11 (cycle == 11);
   //    testOne('b0, 'b010, 'b1000000000000000, 'b01111111111111111111111111111111,
   //            'b01111111111111111111111111111100,
   //            'b00000000000000000000000000000000,
   //            'b01111111111111100000000000000000); //  11: jmp to user mode, PC==0x7FFFFFFC, offset=0x8000
   // endrule
   // rule t12 (cycle == 12);
   //    testOne('b0, 'b010, 'b1111111111110111, 'b10000111011001010100001100100001,
   //            'b00000111011001010100001100100000,
   //            'b00000111011001010100001100100100,
   //            'b00000111011001010100001100000000); //  12: jmp to super mode?, PC==0x07654320,e offset=-9
   // endrule
   // rule t13 (cycle == 13);
   //    testOne('b0, 'b010, 'b0000000000000000, 'b00000000000000000000000000000100,
   //            'b00000000000000000000000000000100,
   //            'b00000000000000000000000000001000,
   //            'b00000000000000000000000000001000); //  13: jmp, PC==0x0
   // endrule
   // rule t14 (cycle == 14);
   //    testOne('b0, 'b000, 'b0000000000000000, 'b00000000000000000000000000000000,
   //            'b00000000000000000000000000001000,
   //            'b00000000000000000000000000001100,
   //            'b00000000000000000000000000001100); //  14: inc
   // endrule
   // rule t15 (cycle == 15);
   //    testOne('b0, 'b000, 'b0000000000000000, 'b00000000000000000000000000000000,
   //            'b00000000000000000000000000001100,
   //            'b00000000000000000000000000010000,
   //            'b00000000000000000000000000010000); //  15: inc
   // endrule
   // rule t16 (cycle == 16);
   //    testOne('b0, 'b000, 'b0000000000000000, 'b00000000000000000000000000000000,
   //            'b00000000000000000000000000010000,
   //            'b00000000000000000000000000010100,
   //            'b00000000000000000000000000010100); //  16: inc
   // endrule
   // rule t17 (cycle == 17);
   //    testOne('b0, 'b001, 'b0000000000000010, 'b00000000000000000000000011110000,
   //            'b00000000000000000000000000011100,
   //            'b00000000000000000000000000100000,
   //            'b00000000000000000000000000101000); //  17: br, offset=3, PC==0x1C
   // endrule
   // rule t18 (cycle == 18);
   //    testOne('b0, 'b000, 'b0000000000000000, 'b00000000000000000000000000000000,
   //            'b00000000000000000000000000100000,
   //            'b00000000000000000000000000100100,
   //            'b00000000000000000000000000100100); //  18: inc
   // endrule
   // rule t19 (cycle == 19);
   //    testOne('b0, 'b010, 'b0000000000000000, 'b00000000000000000000000000111100,
   //            'b00000000000000000000000000111100,
   //            'b00000000000000000000000001000000,
   //            'b00000000000000000000000001000000); //  19: jmp, PC==0x3C
   // endrule
   // rule t20 (cycle == 20);
   //    testOne('b0, 'b000, 'b0000000000000000, 'b00000000000000000000000000000000,
   //            'b00000000000000000000000001000000,
   //            'b00000000000000000000000001000100,
   //            'b00000000000000000000000001000100); //  20: inc
   // endrule
   // rule t21 (cycle == 21);
   //    testOne('b0, 'b010, 'b0000000000000000, 'b00000000000000000000000001111100,
   //            'b00000000000000000000000001111100,
   //            'b00000000000000000000000010000000,
   //            'b00000000000000000000000010000000); //  21: jmp, PC==0x7C
   // endrule
   // rule t22 (cycle == 22);
   //    testOne('b0, 'b000, 'b0000000000000000, 'b00000000000000000000000000000000,
   //            'b00000000000000000000000010000000,
   //            'b00000000000000000000000010000100,
   //            'b00000000000000000000000010000100); //  22: inc
   // endrule
   // rule t23 (cycle == 23);
   //    testOne('b0, 'b010, 'b0000000000000000, 'b00000000000000001111111111111100,
   //            'b00000000000000001111111111111100,
   //            'b00000000000000010000000000000000,
   //            'b00000000000000010000000000000000); //  23: jmp, PC==0xFFFC
   // endrule
   // rule t24 (cycle == 24);
   //    testOne('b0, 'b000, 'b0000000000000000, 'b00000000000000000000000000000000,
   //            'b00000000000000010000000000000000,
   //            'b00000000000000010000000000000100,
   //            'b00000000000000010000000000000100); //  24: inc
   // endrule
   // rule t25 (cycle == 25);
   //    testOne('b0, 'b010, 'b0000000000000000, 'b00000000111111111111111111111100,
   //            'b00000000111111111111111111111100,
   //            'b00000001000000000000000000000000,
   //            'b00000001000000000000000000000000); //  25: jmp, PC==0xFFFFFC
   // endrule
   // rule t26 (cycle == 26);
   //    testOne('b0, 'b000, 'b0000000000000000, 'b00000000000000000000000000000000,
   //            'b00000001000000000000000000000000,
   //            'b00000001000000000000000000000100,
   //            'b00000001000000000000000000000100); //  26: inc
   // endrule
   // rule t27 (cycle == 27);
   //    testOne('b0, 'b010, 'b0000000000000000, 'b01111111111111111111111111111100,
   //            'b01111111111111111111111111111100,
   //            'b00000000000000000000000000000000,
   //            'b00000000000000000000000000000000); //  27: jmp, PC==0x7FFFFFFC
   // endrule
   // rule t28 (cycle == 28);
   //    testOne('b0, 'b000, 'b1111111111111110, 'b00000000000000000000000000000000,
   //            'b00000000000000000000000000000000,
   //            'b00000000000000000000000000000100,
   //            'b01111111111111111111111111111100); //  28: inc
   // endrule
   // rule done (cycle > 1);
   //    $finish();
   // endrule
   
endmodule
