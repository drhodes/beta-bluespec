../cmp/Cmp.bsv