../shift/Shift.bsv