../arith/Arith.bsv