import Ctl::*;

(* synthesize *)
module mkTbCtl(Empty);
   function testOne (Bit#(6) op, Bit#(1) reset, Bit#(1) irq, Bit#(1) z, 
                     Bit#(6) alufn, Bit#(1) asel, Bit#(1) bsel, Bit#(1) moe, 
                     Bit#(1) mwr, Bit#(3) pcsel, Bit#(1) ra2sel, Bit#(1) wasel, 
                     Bit#(2) wdsel, Bit#(1) werf, Integer testnum) = 
   action
      let got = ctl(op, reset, irq, z);
      if (got.alufn != alufn) $display(testnum, " alufn: FAIL got: %b, exp: %b", got.alufn, alufn);
      if (got.alufn == alufn) $display("PASS");
      if (got.asel != asel) $display(testnum, " asel: FAIL got: %b, exp: %b", got.asel, asel);
      if (got.bsel != bsel) $display(testnum, " bsel: FAIL got: %b, exp: %b", got.bsel, bsel);
      if (got.moe != moe) $display(testnum, " moe: FAIL got: %b, exp: %b", got.moe, moe);
      if (got.mwr != mwr) $display(testnum, " mwr: FAIL got: %b, exp: %b", got.mwr, mwr);
      if (got.pcsel != pcsel) $display(testnum, " pcsel: FAIL got: %b, exp: %b", got.pcsel, pcsel);
      if (got.ra2sel != ra2sel) $display(testnum, " ra2sel: FAIL got: %b, exp: %b", got.ra2sel, ra2sel);
      if (got.wasel != wasel) $display(testnum, " wasel: FAIL got: %b, exp: %b", got.wasel, wasel);
      if (got.wdsel != wdsel) $display(testnum, " wdsel: FAIL got: %b, exp: %b", got.wdsel, wdsel);
      if (got.werf != werf) $display(testnum, " werf: FAIL got: %b, exp: %b", got.werf, werf);
   endaction;
   
   rule testAll;
      testOne('b000000, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 1); // 1: op=0b000000 ???
      testOne('b000000, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 2); // 2: op=0b000000 ???
      testOne('b000000, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 3); // 3: op=0b000000 ???
      testOne('b000000, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 4); // 4: op=0b000000 ???
      testOne('b000000, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 5); // 5: op=0b000000 ???
      testOne('b000000, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 6); // 6: op=0b000000 ???
      testOne('b000000, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 7); // 7: op=0b000000 ???
      testOne('b000000, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 8); // 8: op=0b000000 ???
      testOne('b000001, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 9); // 9: op=0b000001 ???
      testOne('b000001, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 10); // 10: op=0b000001 ???
      testOne('b000001, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 11); // 11: op=0b000001 ???
      testOne('b000001, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 12); // 12: op=0b000001 ???
      testOne('b000001, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 13); // 13: op=0b000001 ???
      testOne('b000001, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 14); // 14: op=0b000001 ???
      testOne('b000001, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 15); // 15: op=0b000001 ???
      testOne('b000001, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 16); // 16: op=0b000001 ???
      testOne('b000010, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 17); // 17: op=0b000010 ???
      testOne('b000010, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 18); // 18: op=0b000010 ???
      testOne('b000010, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 19); // 19: op=0b000010 ???
      testOne('b000010, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 20); // 20: op=0b000010 ???
      testOne('b000010, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 21); // 21: op=0b000010 ???
      testOne('b000010, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 22); // 22: op=0b000010 ???
      testOne('b000010, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 23); // 23: op=0b000010 ???
      testOne('b000010, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 24); // 24: op=0b000010 ???
      testOne('b000011, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 25); // 25: op=0b000011 ???
      testOne('b000011, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 26); // 26: op=0b000011 ???
      testOne('b000011, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 27); // 27: op=0b000011 ???
      testOne('b000011, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 28); // 28: op=0b000011 ???
      testOne('b000011, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 29); // 29: op=0b000011 ???
      testOne('b000011, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 30); // 30: op=0b000011 ???
      testOne('b000011, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 31); // 31: op=0b000011 ???
      testOne('b000011, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 32); // 32: op=0b000011 ???
      testOne('b000100, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 33); // 33: op=0b000100 ???
      testOne('b000100, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 34); // 34: op=0b000100 ???
      testOne('b000100, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 35); // 35: op=0b000100 ???
      testOne('b000100, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 36); // 36: op=0b000100 ???
      testOne('b000100, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 37); // 37: op=0b000100 ???
      testOne('b000100, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 38); // 38: op=0b000100 ???
      testOne('b000100, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 39); // 39: op=0b000100 ???
      testOne('b000100, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 40); // 40: op=0b000100 ???
      testOne('b000101, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 41); // 41: op=0b000101 ???
      testOne('b000101, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 42); // 42: op=0b000101 ???
      testOne('b000101, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 43); // 43: op=0b000101 ???
      testOne('b000101, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 44); // 44: op=0b000101 ???
      testOne('b000101, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 45); // 45: op=0b000101 ???
      testOne('b000101, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 46); // 46: op=0b000101 ???
      testOne('b000101, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 47); // 47: op=0b000101 ???
      testOne('b000101, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 48); // 48: op=0b000101 ???
      testOne('b000110, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 49); // 49: op=0b000110 ???
      testOne('b000110, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 50); // 50: op=0b000110 ???
      testOne('b000110, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 51); // 51: op=0b000110 ???
      testOne('b000110, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 52); // 52: op=0b000110 ???
      testOne('b000110, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 53); // 53: op=0b000110 ???
      testOne('b000110, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 54); // 54: op=0b000110 ???
      testOne('b000110, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 55); // 55: op=0b000110 ???
      testOne('b000110, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 56); // 56: op=0b000110 ???
      testOne('b000111, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 57); // 57: op=0b000111 ???
      testOne('b000111, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 58); // 58: op=0b000111 ???
      testOne('b000111, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 59); // 59: op=0b000111 ???
      testOne('b000111, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 60); // 60: op=0b000111 ???
      testOne('b000111, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 61); // 61: op=0b000111 ???
      testOne('b000111, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 62); // 62: op=0b000111 ???
      testOne('b000111, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 63); // 63: op=0b000111 ???
      testOne('b000111, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 64); // 64: op=0b000111 ???
      testOne('b001000, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 65); // 65: op=0b001000 ???
      testOne('b001000, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 66); // 66: op=0b001000 ???
      testOne('b001000, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 67); // 67: op=0b001000 ???
      testOne('b001000, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 68); // 68: op=0b001000 ???
      testOne('b001000, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 69); // 69: op=0b001000 ???
      testOne('b001000, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 70); // 70: op=0b001000 ???
      testOne('b001000, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 71); // 71: op=0b001000 ???
      testOne('b001000, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 72); // 72: op=0b001000 ???
      testOne('b001001, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 73); // 73: op=0b001001 ???
      testOne('b001001, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 74); // 74: op=0b001001 ???
      testOne('b001001, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 75); // 75: op=0b001001 ???
      testOne('b001001, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 76); // 76: op=0b001001 ???
      testOne('b001001, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 77); // 77: op=0b001001 ???
      testOne('b001001, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 78); // 78: op=0b001001 ???
      testOne('b001001, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 79); // 79: op=0b001001 ???
      testOne('b001001, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 80); // 80: op=0b001001 ???
      testOne('b001010, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 81); // 81: op=0b001010 ???
      testOne('b001010, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 82); // 82: op=0b001010 ???
      testOne('b001010, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 83); // 83: op=0b001010 ???
      testOne('b001010, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 84); // 84: op=0b001010 ???
      testOne('b001010, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 85); // 85: op=0b001010 ???
      testOne('b001010, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 86); // 86: op=0b001010 ???
      testOne('b001010, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 87); // 87: op=0b001010 ???
      testOne('b001010, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 88); // 88: op=0b001010 ???
      testOne('b001011, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 89); // 89: op=0b001011 ???
      testOne('b001011, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 90); // 90: op=0b001011 ???
      testOne('b001011, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 91); // 91: op=0b001011 ???
      testOne('b001011, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 92); // 92: op=0b001011 ???
      testOne('b001011, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 93); // 93: op=0b001011 ???
      testOne('b001011, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 94); // 94: op=0b001011 ???
      testOne('b001011, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 95); // 95: op=0b001011 ???
      testOne('b001011, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 96); // 96: op=0b001011 ???
      testOne('b001100, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 97); // 97: op=0b001100 ???
      testOne('b001100, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 98); // 98: op=0b001100 ???
      testOne('b001100, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 99); // 99: op=0b001100 ???
      testOne('b001100, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 100); // 100: op=0b001100 ???
      testOne('b001100, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 101); // 101: op=0b001100 ???
      testOne('b001100, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 102); // 102: op=0b001100 ???
      testOne('b001100, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 103); // 103: op=0b001100 ???
      testOne('b001100, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 104); // 104: op=0b001100 ???
      testOne('b001101, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 105); // 105: op=0b001101 ???
      testOne('b001101, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 106); // 106: op=0b001101 ???
      testOne('b001101, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 107); // 107: op=0b001101 ???
      testOne('b001101, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 108); // 108: op=0b001101 ???
      testOne('b001101, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 109); // 109: op=0b001101 ???
      testOne('b001101, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 110); // 110: op=0b001101 ???
      testOne('b001101, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 111); // 111: op=0b001101 ???
      testOne('b001101, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 112); // 112: op=0b001101 ???
      testOne('b001110, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 113); // 113: op=0b001110 ???
      testOne('b001110, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 114); // 114: op=0b001110 ???
      testOne('b001110, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 115); // 115: op=0b001110 ???
      testOne('b001110, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 116); // 116: op=0b001110 ???
      testOne('b001110, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 117); // 117: op=0b001110 ???
      testOne('b001110, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 118); // 118: op=0b001110 ???
      testOne('b001110, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 119); // 119: op=0b001110 ???
      testOne('b001110, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 120); // 120: op=0b001110 ???
      testOne('b001111, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 121); // 121: op=0b001111 ???
      testOne('b001111, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 122); // 122: op=0b001111 ???
      testOne('b001111, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 123); // 123: op=0b001111 ???
      testOne('b001111, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 124); // 124: op=0b001111 ???
      testOne('b001111, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 125); // 125: op=0b001111 ???
      testOne('b001111, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 126); // 126: op=0b001111 ???
      testOne('b001111, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 127); // 127: op=0b001111 ???
      testOne('b001111, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 128); // 128: op=0b001111 ???
      testOne('b010000, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 129); // 129: op=0b010000 ???
      testOne('b010000, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 130); // 130: op=0b010000 ???
      testOne('b010000, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 131); // 131: op=0b010000 ???
      testOne('b010000, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 132); // 132: op=0b010000 ???
      testOne('b010000, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 133); // 133: op=0b010000 ???
      testOne('b010000, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 134); // 134: op=0b010000 ???
      testOne('b010000, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 135); // 135: op=0b010000 ???
      testOne('b010000, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 136); // 136: op=0b010000 ???
      testOne('b010001, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 137); // 137: op=0b010001 ???
      testOne('b010001, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 138); // 138: op=0b010001 ???
      testOne('b010001, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 139); // 139: op=0b010001 ???
      testOne('b010001, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 140); // 140: op=0b010001 ???
      testOne('b010001, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 141); // 141: op=0b010001 ???
      testOne('b010001, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 142); // 142: op=0b010001 ???
      testOne('b010001, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 143); // 143: op=0b010001 ???
      testOne('b010001, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 144); // 144: op=0b010001 ???
      testOne('b010010, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 145); // 145: op=0b010010 ???
      testOne('b010010, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 146); // 146: op=0b010010 ???
      testOne('b010010, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 147); // 147: op=0b010010 ???
      testOne('b010010, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 148); // 148: op=0b010010 ???
      testOne('b010010, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 149); // 149: op=0b010010 ???
      testOne('b010010, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 150); // 150: op=0b010010 ???
      testOne('b010010, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 151); // 151: op=0b010010 ???
      testOne('b010010, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 152); // 152: op=0b010010 ???
      testOne('b010011, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 153); // 153: op=0b010011 ???
      testOne('b010011, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 154); // 154: op=0b010011 ???
      testOne('b010011, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 155); // 155: op=0b010011 ???
      testOne('b010011, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 156); // 156: op=0b010011 ???
      testOne('b010011, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 157); // 157: op=0b010011 ???
      testOne('b010011, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 158); // 158: op=0b010011 ???
      testOne('b010011, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 159); // 159: op=0b010011 ???
      testOne('b010011, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 160); // 160: op=0b010011 ???
      testOne('b010100, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 161); // 161: op=0b010100 ???
      testOne('b010100, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 162); // 162: op=0b010100 ???
      testOne('b010100, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 163); // 163: op=0b010100 ???
      testOne('b010100, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 164); // 164: op=0b010100 ???
      testOne('b010100, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 165); // 165: op=0b010100 ???
      testOne('b010100, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 166); // 166: op=0b010100 ???
      testOne('b010100, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 167); // 167: op=0b010100 ???
      testOne('b010100, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 168); // 168: op=0b010100 ???
      testOne('b010101, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 169); // 169: op=0b010101 ???
      testOne('b010101, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 170); // 170: op=0b010101 ???
      testOne('b010101, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 171); // 171: op=0b010101 ???
      testOne('b010101, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 172); // 172: op=0b010101 ???
      testOne('b010101, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 173); // 173: op=0b010101 ???
      testOne('b010101, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 174); // 174: op=0b010101 ???
      testOne('b010101, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 175); // 175: op=0b010101 ???
      testOne('b010101, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 176); // 176: op=0b010101 ???
      testOne('b010110, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 177); // 177: op=0b010110 ???
      testOne('b010110, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 178); // 178: op=0b010110 ???
      testOne('b010110, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 179); // 179: op=0b010110 ???
      testOne('b010110, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 180); // 180: op=0b010110 ???
      testOne('b010110, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 181); // 181: op=0b010110 ???
      testOne('b010110, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 182); // 182: op=0b010110 ???
      testOne('b010110, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 183); // 183: op=0b010110 ???
      testOne('b010110, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 184); // 184: op=0b010110 ???
      testOne('b010111, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 185); // 185: op=0b010111 ???
      testOne('b010111, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 186); // 186: op=0b010111 ???
      testOne('b010111, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 187); // 187: op=0b010111 ???
      testOne('b010111, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 188); // 188: op=0b010111 ???
      testOne('b010111, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 189); // 189: op=0b010111 ???
      testOne('b010111, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 190); // 190: op=0b010111 ???
      testOne('b010111, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 191); // 191: op=0b010111 ???
      testOne('b010111, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 192); // 192: op=0b010111 ???
      testOne('b011000, 0,0,0, 'b010000, 0, 1, 1, 0, 'b000, ?, 0, 'b10, 1, 193); // 193: op=0b011000 0D
      testOne('b011000, 0,0,1, 'b010000, 0, 1, 1, 0, 'b000, ?, 0, 'b10, 1, 194); // 194: op=0b011000 0D
      testOne('b011000, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 195); // 195: op=0b011000 0D
      testOne('b011000, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 196); // 196: op=0b011000 0D
      testOne('b011000, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 197); // 197
      testOne('b011000, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 198); // 198
      testOne('b011000, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 199); // 199
      testOne('b011000, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 200); // 200
      testOne('b011001, 0,0,0, 'b010000, 0, 1, 0, 1, 'b000, 1, ?, ?, 0, 201); // 201
      testOne('b011001, 0,0,1, 'b010000, 0, 1, 0, 1, 'b000, 1, ?, ?, 0, 202); // 202
      testOne('b011001, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 203); // 203
      testOne('b011001, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 204); // 204
      testOne('b011001, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 205); // 205
      testOne('b011001, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 206); // 206
      testOne('b011001, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 207); // 207
      testOne('b011001, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 208); // 208
      testOne('b011010, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 209); // 209
      testOne('b011010, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 210); // 210
      testOne('b011010, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 211); // 211
      testOne('b011010, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 212); // 212
      testOne('b011010, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 213); // 213
      testOne('b011010, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 214); // 214
      testOne('b011010, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 215); // 215
      testOne('b011010, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 216); // 216
      testOne('b011011, 0,0,0, ?, ?, ?, ?, 0, 'b010, ?, 0, 'b00, 1, 217); // 217
      testOne('b011011, 0,0,1, ?, ?, ?, ?, 0, 'b010, ?, 0, 'b00, 1, 218); // 218
      testOne('b011011, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 219); // 219
      testOne('b011011, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 220); // 220
      testOne('b011011, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 221); // 221
      testOne('b011011, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 222); // 222
      testOne('b011011, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 223); // 223
      testOne('b011011, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 224); // 224
      testOne('b011100, 0,0,0, ?, ?, ?, ?, 0, 'b000, ?, 0, 'b00, 1, 225); // 225
      testOne('b011100, 0,0,1, ?, ?, ?, ?, 0, 'b001, ?, 0, 'b00, 1, 226); // 226
      testOne('b011100, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 227); // 227
      testOne('b011100, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 228); // 228
      testOne('b011100, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 229); // 229
      testOne('b011100, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 230); // 230
      testOne('b011100, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 231); // 231
      testOne('b011100, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 232); // 232
      testOne('b011101, 0,0,0, ?, ?, ?, ?, 0, 'b001, ?, 0, 'b00, 1, 233); // 233
      testOne('b011101, 0,0,1, ?, ?, ?, ?, 0, 'b000, ?, 0, 'b00, 1, 234); // 234
      testOne('b011101, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 235); // 235
      testOne('b011101, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 236); // 236
      testOne('b011101, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 237); // 237
      testOne('b011101, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 238); // 238
      testOne('b011101, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 239); // 239
      testOne('b011101, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 240); // 240
      testOne('b011110, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 241); // 241
      testOne('b011110, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 242); // 242
      testOne('b011110, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 243); // 243
      testOne('b011110, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 244); // 244
      testOne('b011110, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 245); // 245
      testOne('b011110, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 246); // 246
      testOne('b011110, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 247); // 247
      testOne('b011110, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 248); // 248
      testOne('b011111, 0,0,0, 'b101010, 1, ?, 1, 0, 'b000, ?, 0, 'b10, 1, 249); // 249
      testOne('b011111, 0,0,1, 'b101010, 1, ?, 1, 0, 'b000, ?, 0, 'b10, 1, 250); // 250
      testOne('b011111, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 251); // 251
      testOne('b011111, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 252); // 252
      testOne('b011111, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 253); // 253
      testOne('b011111, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 254); // 254
      testOne('b011111, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 255); // 255
      testOne('b011111, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 256); // 256
      testOne('b100000, 0,0,0, 'b010000, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 257); // 257
      testOne('b100000, 0,0,1, 'b010000, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 258); // 258
      testOne('b100000, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 259); // 259
      testOne('b100000, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 260); // 260
      testOne('b100000, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 261); // 261
      testOne('b100000, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 262); // 262
      testOne('b100000, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 263); // 263
      testOne('b100000, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 264); // 264
      testOne('b100001, 0,0,0, 'b010001, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 265); // 265
      testOne('b100001, 0,0,1, 'b010001, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 266); // 266
      testOne('b100001, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 267); // 267
      testOne('b100001, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 268); // 268
      testOne('b100001, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 269); // 269
      testOne('b100001, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 270); // 270
      testOne('b100001, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 271); // 271
      testOne('b100001, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 272); // 272
      testOne('b100010, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 273); // 273
      testOne('b100010, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 274); // 274
      testOne('b100010, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 275); // 275
      testOne('b100010, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 276); // 276
      testOne('b100010, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 277); // 277
      testOne('b100010, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 278); // 278
      testOne('b100010, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 279); // 279
      testOne('b100010, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 280); // 280
      testOne('b100011, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 281); // 281
      testOne('b100011, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 282); // 282
      testOne('b100011, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 283); // 283
      testOne('b100011, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 284); // 284
      testOne('b100011, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 285); // 285
      testOne('b100011, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 286); // 286
      testOne('b100011, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 287); // 287
      testOne('b100011, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 288); // 288
      testOne('b100100, 0,0,0, 'b000011, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 289); // 289
      testOne('b100100, 0,0,1, 'b000011, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 290); // 290
      testOne('b100100, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 291); // 291
      testOne('b100100, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 292); // 292
      testOne('b100100, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 293); // 293
      testOne('b100100, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 294); // 294
      testOne('b100100, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 295); // 295
      testOne('b100100, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 296); // 296
      testOne('b100101, 0,0,0, 'b000101, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 297); // 297
      testOne('b100101, 0,0,1, 'b000101, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 298); // 298
      testOne('b100101, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 299); // 299
      testOne('b100101, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 300); // 300
      testOne('b100101, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 301); // 301
      testOne('b100101, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 302); // 302
      testOne('b100101, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 303); // 303
      testOne('b100101, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 304); // 304
      testOne('b100110, 0,0,0, 'b000111, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 305); // 305
      testOne('b100110, 0,0,1, 'b000111, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 306); // 306
      testOne('b100110, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 307); // 307
      testOne('b100110, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 308); // 308
      testOne('b100110, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 309); // 309
      testOne('b100110, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 310); // 310
      testOne('b100110, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 311); // 311
      testOne('b100110, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 312); // 312
      testOne('b100111, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 313); // 313
      testOne('b100111, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 314); // 314
      testOne('b100111, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 315); // 315
      testOne('b100111, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 316); // 316
      testOne('b100111, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 317); // 317
      testOne('b100111, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 318); // 318
      testOne('b100111, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 319); // 319
      testOne('b100111, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 320); // 320
      testOne('b101000, 0,0,0, 'b101000, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 321); // 321
      testOne('b101000, 0,0,1, 'b101000, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 322); // 322
      testOne('b101000, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 323); // 323
      testOne('b101000, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 324); // 324
      testOne('b101000, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 325); // 325
      testOne('b101000, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 326); // 326
      testOne('b101000, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 327); // 327
      testOne('b101000, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 328); // 328
      testOne('b101001, 0,0,0, 'b101110, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 329); // 329
      testOne('b101001, 0,0,1, 'b101110, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 330); // 330
      testOne('b101001, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 331); // 331
      testOne('b101001, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 332); // 332
      testOne('b101001, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 333); // 333
      testOne('b101001, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 334); // 334
      testOne('b101001, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 335); // 335
      testOne('b101001, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 336); // 336
      testOne('b101010, 0,0,0, 'b100110, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 337); // 337
      testOne('b101010, 0,0,1, 'b100110, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 338); // 338
      testOne('b101010, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 339); // 339
      testOne('b101010, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 340); // 340
      testOne('b101010, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 341); // 341
      testOne('b101010, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 342); // 342
      testOne('b101010, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 343); // 343
      testOne('b101010, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 344); // 344
      testOne('b101011, 0,0,0, 'b101001, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 345); // 345
      testOne('b101011, 0,0,1, 'b101001, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 346); // 346
      testOne('b101011, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 347); // 347
      testOne('b101011, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 348); // 348
      testOne('b101011, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 349); // 349
      testOne('b101011, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 350); // 350
      testOne('b101011, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 351); // 351
      testOne('b101011, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 352); // 352
      testOne('b101100, 0,0,0, 'b110000, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 353); // 353
      testOne('b101100, 0,0,1, 'b110000, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 354); // 354
      testOne('b101100, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 355); // 355
      testOne('b101100, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 356); // 356
      testOne('b101100, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 357); // 357
      testOne('b101100, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 358); // 358
      testOne('b101100, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 359); // 359
      testOne('b101100, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 360); // 360
      testOne('b101101, 0,0,0, 'b110001, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 361); // 361
      testOne('b101101, 0,0,1, 'b110001, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 362); // 362
      testOne('b101101, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 363); // 363
      testOne('b101101, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 364); // 364
      testOne('b101101, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 365); // 365
      testOne('b101101, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 366); // 366
      testOne('b101101, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 367); // 367
      testOne('b101101, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 368); // 368
      testOne('b101110, 0,0,0, 'b110011, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 369); // 369
      testOne('b101110, 0,0,1, 'b110011, 0, 0, ?, 0, 'b000, 0, 0, 'b01, 1, 370); // 370
      testOne('b101110, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 371); // 371
      testOne('b101110, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 372); // 372
      testOne('b101110, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 373); // 373
      testOne('b101110, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 374); // 374
      testOne('b101110, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 375); // 375
      testOne('b101110, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 376); // 376
      testOne('b101111, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 377); // 377
      testOne('b101111, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 378); // 378
      testOne('b101111, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 379); // 379
      testOne('b101111, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 380); // 380
      testOne('b101111, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 381); // 381
      testOne('b101111, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 382); // 382
      testOne('b101111, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 383); // 383
      testOne('b101111, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 384); // 384
      testOne('b110000, 0,0,0, 'b010000, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 385); // 385
      testOne('b110000, 0,0,1, 'b010000, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 386); // 386
      testOne('b110000, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 387); // 387
      testOne('b110000, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 388); // 388
      testOne('b110000, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 389); // 389
      testOne('b110000, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 390); // 390
      testOne('b110000, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 391); // 391
      testOne('b110000, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 392); // 392
      testOne('b110001, 0,0,0, 'b010001, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 393); // 393
      testOne('b110001, 0,0,1, 'b010001, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 394); // 394
      testOne('b110001, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 395); // 395
      testOne('b110001, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 396); // 396
      testOne('b110001, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 397); // 397
      testOne('b110001, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 398); // 398
      testOne('b110001, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 399); // 399
      testOne('b110001, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 400); // 400
      testOne('b110010, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 401); // 401
      testOne('b110010, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 402); // 402
      testOne('b110010, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 403); // 403
      testOne('b110010, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 404); // 404
      testOne('b110010, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 405); // 405
      testOne('b110010, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 406); // 406
      testOne('b110010, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 407); // 407
      testOne('b110010, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 408); // 408
      testOne('b110011, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 409); // 409
      testOne('b110011, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 410); // 410
      testOne('b110011, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 411); // 411
      testOne('b110011, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 412); // 412
      testOne('b110011, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 413); // 413
      testOne('b110011, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 414); // 414
      testOne('b110011, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 415); // 415
      testOne('b110011, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 416); // 416
      testOne('b110100, 0,0,0, 'b000011, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 417); // 417
      testOne('b110100, 0,0,1, 'b000011, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 418); // 418
      testOne('b110100, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 419); // 419
      testOne('b110100, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 420); // 420
      testOne('b110100, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 421); // 421
      testOne('b110100, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 422); // 422
      testOne('b110100, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 423); // 423
      testOne('b110100, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 424); // 424
      testOne('b110101, 0,0,0, 'b000101, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 425); // 425
      testOne('b110101, 0,0,1, 'b000101, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 426); // 426
      testOne('b110101, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 427); // 427
      testOne('b110101, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 428); // 428
      testOne('b110101, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 429); // 429
      testOne('b110101, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 430); // 430
      testOne('b110101, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 431); // 431
      testOne('b110101, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 432); // 432
      testOne('b110110, 0,0,0, 'b000111, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 433); // 433
      testOne('b110110, 0,0,1, 'b000111, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 434); // 434
      testOne('b110110, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 435); // 435
      testOne('b110110, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 436); // 436
      testOne('b110110, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 437); // 437
      testOne('b110110, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 438); // 438
      testOne('b110110, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 439); // 439
      testOne('b110110, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 440); // 440
      testOne('b110111, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 441); // 441
      testOne('b110111, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 442); // 442
      testOne('b110111, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 443); // 443
      testOne('b110111, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 444); // 444
      testOne('b110111, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 445); // 445
      testOne('b110111, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 446); // 446
      testOne('b110111, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 447); // 447
      testOne('b110111, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 448); // 448
      testOne('b111000, 0,0,0, 'b101000, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 449); // 449
      testOne('b111000, 0,0,1, 'b101000, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 450); // 450
      testOne('b111000, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 451); // 451
      testOne('b111000, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 452); // 452
      testOne('b111000, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 453); // 453
      testOne('b111000, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 454); // 454
      testOne('b111000, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 455); // 455
      testOne('b111000, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 456); // 456
      testOne('b111001, 0,0,0, 'b101110, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 457); // 457
      testOne('b111001, 0,0,1, 'b101110, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 458); // 458
      testOne('b111001, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 459); // 459
      testOne('b111001, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 460); // 460
      testOne('b111001, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 461); // 461
      testOne('b111001, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 462); // 462
      testOne('b111001, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 463); // 463
      testOne('b111001, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 464); // 464
      testOne('b111010, 0,0,0, 'b100110, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 465); // 465
      testOne('b111010, 0,0,1, 'b100110, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 466); // 466
      testOne('b111010, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 467); // 467
      testOne('b111010, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 468); // 468
      testOne('b111010, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 469); // 469
      testOne('b111010, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 470); // 470
      testOne('b111010, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 471); // 471
      testOne('b111010, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 472); // 472
      testOne('b111011, 0,0,0, 'b101001, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 473); // 473
      testOne('b111011, 0,0,1, 'b101001, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 474); // 474
      testOne('b111011, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 475); // 475
      testOne('b111011, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 476); // 476
      testOne('b111011, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 477); // 477
      testOne('b111011, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 478); // 478
      testOne('b111011, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 479); // 479
      testOne('b111011, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 480); // 480
      testOne('b111100, 0,0,0, 'b110000, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 481); // 481
      testOne('b111100, 0,0,1, 'b110000, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 482); // 482
      testOne('b111100, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 483); // 483
      testOne('b111100, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 484); // 484
      testOne('b111100, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 485); // 485
      testOne('b111100, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 486); // 486
      testOne('b111100, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 487); // 487
      testOne('b111100, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 488); // 488
      testOne('b111101, 0,0,0, 'b110001, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 489); // 489
      testOne('b111101, 0,0,1, 'b110001, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 490); // 490
      testOne('b111101, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 491); // 491
      testOne('b111101, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 492); // 492
      testOne('b111101, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 493); // 493
      testOne('b111101, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 494); // 494
      testOne('b111101, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 495); // 495
      testOne('b111101, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 496); // 496
      testOne('b111110, 0,0,0, 'b110011, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 497); // 497
      testOne('b111110, 0,0,1, 'b110011, 0, 1, ?, 0, 'b000, ?, 0, 'b01, 1, 498); // 498
      testOne('b111110, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 499); // 499
      testOne('b111110, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 500); // 500
      testOne('b111110, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 501); // 501
      testOne('b111110, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 502); // 502
      testOne('b111110, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 503); // 503
      testOne('b111110, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 504); // 504
      testOne('b111111, 0,0,0, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 505); // 505
      testOne('b111111, 0,0,1, ?, ?, ?, ?, 0, 'b011, ?, 1, 'b00, 1, 506); // 506
      testOne('b111111, 0,1,0, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 507); // 507
      testOne('b111111, 0,1,1, ?, ?, ?, ?, 0, 'b100, ?, 1, 'b00, 1, 508); // 508
      testOne('b111111, 1,0,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 509); // 509
      testOne('b111111, 1,0,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 510); // 510
      testOne('b111111, 1,1,0, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 511); // 511
      testOne('b111111, 1,1,1, ?, ?, ?, ?, 0, ?, ?, ?, ?, ?, 512); // 512
      
      $finish();
   endrule
endmodule
