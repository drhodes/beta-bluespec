../bool/Bool.bsv