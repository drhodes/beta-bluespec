import Memory::*;
import BRAMFIFO::*;

typedef struct {
   Bit#(6) alufn;
   Bit#(1) asel;
   Bit#(1) bsel;
   Bit#(1) moe;
   Bit#(1) mwr;
   Bit#(3) pcsel;
   Bit#(1) ra2sel;
   Bit#(1) wasel;
   Bit#(2) wdsel;
   Bit#(1) werf;
} CtlOut deriving (Bits, Eq, FShow);


function CtlOut g (Bit#(18) xs);
   return CtlOut{alufn:xs[17:12], asel:xs[11], bsel:xs[10], moe:xs[9], mwr:xs[8], 
            pcsel:xs[7:5], ra2sel:xs[4], wasel:xs[3], wdsel:xs[2:1], werf:xs[0]};
endfunction

function CtlOut ctl (Bit#(6) op, Bit#(1) reset, Bit#(1) irq, Bit#(1) z);
   let out = case (op)
      //            alufn[17:12]
      //            |     asel, bsel
      //            |     | moe, mwr
      //            |     | | pcsel[2:0]
      //            |     | | |  ra2sel
      //            |     | | |  | wasel, wdsel[1:0], werf
      //            |     | | |  | |
      'b000000: g('b000000000001101001);  // 
      'b000001: g('b000000000001101001);  // 
      'b000010: g('b000000000001101001);  // 
      'b000011: g('b000000000001101001);  // 
      'b000100: g('b000000000001101001);  // 
      'b000101: g('b000000000001101001);  // 
      'b000110: g('b000000000001101001);  // 
      'b000111: g('b000000000001101001);  // 
      'b001000: g('b000000000001101001);  // 
      'b001001: g('b000000000001101001);  // 
      'b001010: g('b000000000001101001);  // 
      'b001011: g('b000000000001101001);  // 
      'b001100: g('b000000000001101001);  // 
      'b001101: g('b000000000001101001);  // 
      'b001110: g('b000000000001101001);  // 
      'b001111: g('b000000000001101001);  // 
      'b010000: g('b000000000001101001);  // 
      'b010001: g('b000000000001101001);  // 
      'b010010: g('b000000000001101001);  // 
      'b010011: g('b000000000001101001);  // 
      'b010100: g('b000000000001101001);  // 
      'b010101: g('b000000000001101001);  // 
      'b010110: g('b000000000001101001);  // 
      'b010111: g('b000000000001101001);  // 
      'b011000: g('b010000011000000101);  // 
      'b011001: g('b010000010100010000);  // ST *
      'b011010: g('b000000000001101001);  
      'b011011: g('b000000000001000001); // JMP *
      'b011100: g('b000000000000000001); // BEQ, Z01:0, submod handles pcsel *
      'b011101: g('b000000000000000001); // BNE, Z00:1, submod handles pcsel *
      'b011110: g('b000000000001101001); 
      'b011111: g('b101010101000000101); // LDR *
      'b100000: g('b010000000000000011); // ADD
      'b100001: g('b010001000000000011); // SUB
      'b100010: g('b000000000001101001); // [normally MUL, but ILLOP for our ALU]
      'b100011: g('b000000000001101001); // [normally DIV, but ILOOP for our ALU]
      'b100100: g('b000011000000000011); // CMPEQ
      'b100101: g('b000101000000000011); // CMPLT
      'b100110: g('b000111000000000011); // CMPLE
      'b100111: g('b000000000001101001); 
      'b101000: g('b101000000000000011); // AND
      'b101001: g('b101110000000000011); // OR
      'b101010: g('b100110000000000011); // XOR
      'b101011: g('b101001000000000011); // XNOR
      'b101100: g('b110000000000000011); // SHL
      'b101101: g('b110001000000000011); // SHR
      'b101110: g('b110011000000000011); // SRA
      'b101111: g('b000000000001101001);  
      'b110000: g('b010000010000000011); // ADDC
      'b110001: g('b010001010000000011); // SUBC
      'b110010: g('b000000000001101001); // [normally MULC, but ILLOP for our ALU]
      'b110011: g('b000000000001101001); // [normally DIVC, but ILLOP for our ALU]
      'b110100: g('b000011010000000011); // CMPEQC
      'b110101: g('b000101010000000011); // CMPLTC
      'b110110: g('b000111010000000011); // CMPLEC
      'b110111: g('b000000000001101001); //  
      'b111000: g('b101000010000000011); // ANDC
      'b111001: g('b101110010000000011); // ORC
      'b111010: g('b100110010000000011); // XORC
      'b111011: g('b101001010000000011); // XNORC
      'b111100: g('b110000010000000011); // SHLC
      'b111101: g('b110001010000000011); // SHRC
      'b111110: g('b110011010000000011); // SRAC
      'b111111: g('b000000000001101001); //  
   endcase;

   
   //$display("ASDF", out);
   
   if (irq == 1) begin
      out.werf = 1;
      out.wasel = 1;
      out.wdsel = 'b00;
      out.pcsel = 'b100;
   end
   
   if (reset == 1) out.mwr = 0;
   else if (reset == 0 && irq == 1) out.mwr = 0;
   
   let br_beq = ~op[5] & op[4] & op[3] & op[2] & ~op[1] & ~op[0];
   let br_bne = ~op[5] & op[4] & op[3] & op[2] & ~op[1] & op[0];
   
   let is_branch_instr = br_beq | br_bne;
   let br_taken = (z & br_beq) | (~z & br_bne);

   if (irq == 0 && is_branch_instr == 1) begin
      if (br_taken == 1) out.pcsel = 'b001;
      else out.pcsel = 'b000;
   end
      
   
   
   
   return out;
endfunction
      // //                   alufn[17:12]
      // //                   |     asel, bsel
      // //                   |     | moe, mwr
      // //                   |     | | pcsel[2:0]
      // //                   |     | | |  ra2sel
      // //                   |     | | |  | wasel, wdsel[1:0], werf
      // //                   |     | | |  | |
      // 'b000000: return g('b?????????0011?1001);  // 
      // 'b000001: return g('b?????????0011?1001);  // 
      // 'b000010: return g('b?????????0011?1001);  // 
      // 'b000011: return g('b?????????0011?1001);  // 
      // 'b000100: return g('b?????????0011?1001);  // 
      // 'b000101: return g('b?????????0011?1001);  // 
      // 'b000110: return g('b?????????0011?1001);  // 
      // 'b000111: return g('b?????????0011?1001);  // 
      // 'b001000: return g('b?????????0011?1001);  // 
      // 'b001001: return g('b?????????0011?1001);  // 
      // 'b001010: return g('b?????????0011?1001);  // 
      // 'b001011: return g('b?????????0011?1001);  // 
      // 'b001100: return g('b?????????0011?1001);  // 
      // 'b001101: return g('b?????????0011?1001);  // 
      // 'b001110: return g('b?????????0011?1001);  // 
      // 'b001111: return g('b?????????0011?1001);  // 
      // 'b010000: return g('b?????????0011?1001);  // 
      // 'b010001: return g('b?????????0011?1001);  // 
      // 'b010010: return g('b?????????0011?1001);  // 
      // 'b010011: return g('b?????????0011?1001);  // 
      // 'b010100: return g('b?????????0011?1001);  // 
      // 'b010101: return g('b?????????0011?1001);  // 
      // 'b010110: return g('b?????????0011?1001);  // 
      // 'b010111: return g('b?????????0011?1001);  // 
      // 'b011000: return g('b0100000110000?0101);  // 
      // 'b011001: return g('b01000001010001???0);  // ST *
      // 'b011010: return g('b?????????0011?1001);  
      // 'b011011: return g('b?????????0010?0001);  // JMP *
      // 'b011100: return g('b?????????0????0001);   //BEQ, Z?1:0, submod handles pcsel *
      // 'b011101: return g('b?????????0????0001);   //BNE, Z?0:1, submod handles pcsel *
      // 'b011110: return g('b?????????0011?1001);  
      // 'b011111: return g('b1010101?10000?0101);   //LDR *
      // 'b100000: return g('b010000000000000011);   //ADD
      // 'b100001: return g('b010001000000000011);   //SUB
      // 'b100010: return g('b?????????0011?1001);   //[normally MUL, but ILLOP for our ALU]
      // 'b100011: return g('b?????????0011?1001);   //[normally DIV, but ILOOP for our ALU]
      // 'b100100: return g('b000011000000000011); //CMPEQ
      // 'b100101: return g('b000101000000000011); //CMPLT
      // 'b100110: return g('b000111000000000011); //CMPLE
      // 'b100111: return g('b?????????0011?1001);  
      // 'b101000: return g('b101000000000000011); // AND
      // 'b101001: return g('b101110000000000011); // OR
      // 'b101010: return g('b100110000000000011); //XOR
      // 'b101011: return g('b101001000000000011); //XNOR
      // 'b101100: return g('b110000000000000011); // SHL
      // 'b101101: return g('b110001000000000011); // SHR
      // 'b101110: return g('b110011000000000011); // SRA
      // 'b101111: return g('b?????????0011?1001);  
      // 'b110000: return g('b010000010000000011); // ADDC
      // 'b110001: return g('b010001010000000011); // SUBC
      // 'b110010: return g('b?????????0011?1001); // [normally MULC, but ILLOP for our ALU]
      // 'b110011: return g('b?????????0011?1001); //   [normally DIVC, but ILLOP for our ALU]
      // 'b110100: return g('b000011010000000011); //   CMPEQC
      // 'b110101: return g('b000101010000000011); //   CMPLTC
      // 'b110110: return g('b000111010000000011); //   CMPLEC
      // 'b110111: return g('b?????????0011?1001); //  
      // 'b111000: return g('b101000010000000011); //   ANDC
      // 'b111001: return g('b101110010000000011); //   ORC
      // 'b111010: return g('b100110010000000011); //   XORC
      // 'b111011: return g('b101001010000000011); //   XNORC
      // 'b111100: return g('b110000010000000011); //   SHLC
      // 'b111101: return g('b110001010000000011); //   SHRC
      // 'b111110: return g('b110011010000000011); //   SRAC
      // 'b111111: return g('b?????????0011?1001); //  




// //alufn[17:12]
// //|      asel, bsel
// //|      |  moe, mwr
// //|      |  |  pcsel[2:0]
// //|      |  |  |   ra2sel
// //|      |  |  |   | wasel, wdsel[1:0], werf
// //|      |  |  |   | |
// 0b??????_??_?0_011_?_1001  // 0b000000
// 0b??????_??_?0_011_?_1001  // 0b000001
// 0b??????_??_?0_011_?_1001  // 0b000010
// 0b??????_??_?0_011_?_1001  // 0b000011
// 0b??????_??_?0_011_?_1001  // 0b000100
// 0b??????_??_?0_011_?_1001  // 0b000101 
// 0b??????_??_?0_011_?_1001  // 0b000110
// 0b??????_??_?0_011_?_1001  // 0b000111

// 0b??????_??_?0_011_?_1001  // 0b001000
// 0b??????_??_?0_011_?_1001  // 0b001001
// 0b??????_??_?0_011_?_1001  // 0b001010
// 0b??????_??_?0_011_?_1001  // 0b001011
// 0b??????_??_?0_011_?_1001  // 0b001100
// 0b??????_??_?0_011_?_1001  // 0b001101
// 0b??????_??_?0_011_?_1001  // 0b001110
// 0b??????_??_?0_011_?_1001  // 0b001111

// //alufn[5:0]
// //|      asel, bsel
// //|      |  moe, mwr
// //|      |  |  pcsel[2:0]
// //|      |  |  |   ra2sel
// //|      |  |  |   | wasel, wdsel[1:0], werf
// //|      |  |  |   | |
// 0b??????_??_?0_011_?_1001  // 0b010000
// 0b??????_??_?0_011_?_1001  // 0b010001
// 0b??????_??_?0_011_?_1001  // 0b010010
// 0b??????_??_?0_011_?_1001  // 0b010011
// 0b??????_??_?0_011_?_1001  // 0b010100
// 0b??????_??_?0_011_?_1001  // 0b010101
// 0b??????_??_?0_011_?_1001  // 0b010110
// 0b??????_??_?0_011_?_1001  // 0b010111

// 0b010000_01_10_000_?_0101  // 0b011000 LD *

// 0b010000_01_01_000_1_???0  // 0b011001 ST *
// 0b??????_??_?0_011_?_1001  // 0b011010
// 0b??????_??_?0_010_?_0001  // 0b011011 JMP *

// 0b??????_??_?0_???_?_0001  // 0b011100 BEQ, Z?1:0, submod handles pcsel *
// 0b??????_??_?0_???_?_0001  // 0b011101 BNE, Z?0:1, submod handles pcsel *

// 0b??????_??_?0_011_?_1001  // 0b011110
// 0b101010_1?_10_000_?_0101  // 0b011111 LDR *

// //alufn[5:0]
// //|      asel, bsel
// //|      |  moe, mwr
// //|      |  |  pcsel[2:0]
// //|      |  |  |   ra2sel
// //|      |  |  |   | wasel, wdsel[1:0], werf
// //|      |  |  |   | |
// 0b010000_00_00_000_0_0011  // 0b100000 ADD
// 0b010001_00_00_000_0_0011  // 0b100001 SUB
// 0b??????_??_?0_011_?_1001  // 0b100010 [normally MUL, but ILLOP for our ALU]
// 0b??????_??_?0_011_?_1001  // 0b100011 [normally DIV, but ILOOP for our ALU]
// 0b000011_00_00_000_0_0011  // 0b100100 CMPEQ
// 0b000101_00_00_000_0_0011  // 0b100101 CMPLT
// 0b000111_00_00_000_0_0011  // 0b100110 CMPLE
// 0b??????_??_?0_011_?_1001  // 0b100111

// 0b101000_00_00_000_0_0011  // 0b101000 AND
// 0b101110_00_00_000_0_0011  // 0b101001 OR
// 0b100110_00_00_000_0_0011  // 0b101010 XOR
// 0b101001_00_00_000_0_0011  // 0b101011 XNOR
// 0b110000_00_00_000_0_0011  // 0b101100 SHL
// 0b110001_00_00_000_0_0011  // 0b101101 SHR
// 0b110011_00_00_000_0_0011  // 0b101110 SRA
// 0b??????_??_?0_011_?_1001  // 0b101111

// //alufn[5:0]
// //|      asel, bsel
// //|      |  moe, mwr
// //|      |  |  pcsel[2:0]
// //|      |  |  |   ra2sel
// //|      |  |  |   | wasel, wdsel[1:0], werf
// //|      |  |  |   | |
// 0b010000_01_00_000_0_0011  // 0b110000 ADDC
// 0b010001_01_00_000_0_0011  // 0b110001 SUBC
// 0b??????_??_?0_011_?_1001  // 0b110010 [normally MULC, but ILLOP for our ALU]
// 0b??????_??_?0_011_?_1001  // 0b110011 [normally DIVC, but ILLOP for our ALU]
// 0b000011_01_00_000_0_0011  // 0b110100 CMPEQC
// 0b000101_01_00_000_0_0011  // 0b110101 CMPLTC
// 0b000111_01_00_000_0_0011  // 0b110110 CMPLEC
// 0b??????_??_?0_011_?_1001  // 0b110111

// 0b101000_01_00_000_0_0011  // 0b111000 ANDC
// 0b101110_01_00_000_0_0011  // 0b111001 ORC
// 0b100110_01_00_000_0_0011  // 0b111010 XORC
// 0b101001_01_00_000_0_0011  // 0b111011 XNORC
// 0b110000_01_00_000_0_0011  // 0b111100 SHLC
// 0b110001_01_00_000_0_0011  // 0b111101 SHRC
// 0b110011_01_00_000_0_0011  // 0b111110 SRAC
// 0b??????_??_?0_011_?_1001  // 0b111111
